// Date: YYYY-MM-DD
// Author: Stephen Zhang
// URL: the url to the question

/** Question:
 * <descrpition of question>
 */

module top_module
(
    input logic in,
    output logic out
);

    assign out = ~in;

endmodule

// EOF
